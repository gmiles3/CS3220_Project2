library verilog;
use verilog.vl_types.all;
entity dprf_testbench is
end dprf_testbench;
